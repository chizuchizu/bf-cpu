module matrixLED (
    output wire [7:0] col,
    output wire [2:0] row
);

    assign col = 8'b00000000;
    assign row = 3'b000;

endmodule