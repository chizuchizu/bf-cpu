module main(
    output odata
);

    assign odata = 1'b0;

endmodule