module 74HC04(
    input [5:0] in
    output [5:0] out
)

    assign out = ~in
endmodule